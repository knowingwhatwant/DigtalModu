module QPSK_Mod()